library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity WB is
end WB;

architecture Behavioral of WB is

begin

-- tratar do DA, WE, DATA do register file neste andar

OLA AMIGOSOSOSOSS


end Behavioral;

